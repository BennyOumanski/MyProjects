LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
LIBRARY altera_mf;
USE altera_mf.altera_mf_components.all;

ENTITY Ifetch IS
	GENERIC (MemWidth	: INTEGER;
			 SIM 		: BOOLEAN);
	PORT(	Instruction							   	: OUT	STD_LOGIC_VECTOR( 31 DOWNTO 0 );
        	PC_plus_4_out 						   	: OUT	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
        	Add_result 							   	: IN 	STD_LOGIC_VECTOR( 7 DOWNTO 0 );
        	PCSrc 								   	: IN 	STD_LOGIC_VECTOR( 1 DOWNTO 0 );
      		PC_out 								   	: OUT	STD_LOGIC_VECTOR( 9 DOWNTO 0 );
			JumpAddr							   	: IN	STD_LOGIC_VECTOR( 7 DOWNTO 0 );
        	clock, ena, Stall_IF,  reset 			: IN 	STD_LOGIC;
			INTA									: IN	STD_LOGIC;
			Read_ISR_PC								: IN	STD_LOGIC;
			HOLD_PC									: IN 	STD_LOGIC;
			ISRAddr									: IN	STD_LOGIC_VECTOR(31 DOWNTO 0)
			);
END Ifetch;

ARCHITECTURE behavior OF Ifetch IS
	SIGNAL PC, PC_plus_4 	 : STD_LOGIC_VECTOR( 9 DOWNTO 0 );
	SIGNAL next_PC			 : STD_LOGIC_VECTOR( 7 DOWNTO 0 );
	SIGNAL Mem_Addr 		 : STD_LOGIC_VECTOR( MemWidth-1 DOWNTO 0 );
	SIGNAL Mem_clock		 : STD_LOGIC;
BEGIN

inst_memory: altsyncram
	
	GENERIC MAP (
		operation_mode => "ROM",
		width_a => 32,
		widthad_a => MemWidth,
		lpm_type => "altsyncram",
		numwords_a             => 2**MemWidth, 
		outdata_reg_a => "UNREGISTERED",
		init_file => "C:\Benny\VHDL\Final Project\Our Project\DataFiles\ITCM.hex",
		intended_device_family => "Cyclone",
		ram_block_type        => "M9K",
		lpm_hint              => "ENABLE_RUNTIME_MOD=YES, INSTANCE_NAME=ITCM"
	)
	PORT MAP (
		clock0     => Mem_clock,  -- Falling Edge
		address_a 	=> Mem_Addr, 
		q_a 			=> Instruction
		);

			
		Mem_clock <= not clock;

		PC(1 DOWNTO 0) <= "00";

		PC_out 			<= PC;
		PC_plus_4_out 	<= PC_plus_4;

		
		ModelSim: 
		IF (SIM = TRUE) GENERATE
			Mem_Addr <= "00" & PC(9 downto 2);
		END GENERATE ModelSim;
		
		FPGA: 
		IF (SIM = FALSE) GENERATE
				Mem_Addr <= PC;
		END GENERATE FPGA;
		

		PC_plus_4( 9 DOWNTO 2 )  <= PC( 9 DOWNTO 2 ) + 1;
       	PC_plus_4( 1 DOWNTO 0 )  <= "00";
		

		Next_PC  <= X"00" 				WHEN Reset = '1' 		ELSE
					ISRAddr(9 DOWNTO 2)	WHEN Read_ISR_PC = '1'	ELSE	-- Interrupt!
					Add_result 			WHEN PCSrc = "01" 		ELSE 	-- branch
					JumpAddr			WHEN PCSrc = "10"		ELSE	-- jump
					PC_plus_4(9 DOWNTO 2);
			

					PROCESS  BEGIN
		WAIT UNTIL ( clock'EVENT ) AND ( clock = '1' );
		IF reset = '1' THEN
			   PC( 9 DOWNTO 2) <= "00000000"; 
		ELSIF (ena = '1' AND Stall_IF = '0' AND HOLD_PC = '0') THEN
			   PC( 9 DOWNTO 2 ) <= next_PC;
		END IF;
	END PROCESS;
END behavior;


